module test(
    a,b,c
);
    input a;
    input b;
    output reg c;
    always @(*) begin
        c = a * b;
        
    end
endmodule

����ļ�һ��lint���