
module if (
    input                 clk     ,
    input                 rst     ,
    input      [31:0]     inst    ,
    input                 jr      ,
    input      [31:0]     jpc     ,
    input                 bhazard ,
    input      [31:0]     bpc     ,
    output     [31:0]     pc      ,
    output     [31:0]     if_inst
);


    
    
endmodule